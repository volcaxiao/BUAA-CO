`timescale 1ns / 1ps

////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer:
//
// Create Date:   17:00:53 10/10/2022
// Design Name:   BlockChecker
// Module Name:   /media/shared/p1/6_BlockChecker/BlockChecker/BlockCheck_tb.v
// Project Name:  BlockChecker
// Target Device:  
// Tool versions:  
// Description: 
//
// Verilog Test Fixture created by ISE for module: BlockChecker
//
// Dependencies:
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
////////////////////////////////////////////////////////////////////////////////

module BlockCheck_tb;

	// Inputs
	reg clk;
	reg reset;
	reg [7:0] in;

	// Outputs
	wire result;

	// Instantiate the Unit Under Test (UUT)
	BlockChecker uut (
		.clk        (clk), 
		.reset      (reset), 
		.in         (in), 
		.result     (result)
	);

	initial begin
		// Initialize Inputs
		clk = 0;
		reset = 0;
		in = "a";

		// Add stimulus here
        #15 in = " ";
        #10 in = "B";
        #10 in = "E";
        #10 in = "g";
        #10 in = "I";
        #10 in = "n";
        #10 in = " ";
        #10 in = "E";
        #10 in = "n";
        #10 in = "d";
        #10 in = "c";
        #10 in = " ";
        #10 in = "e";
        #10 in = "n";
        #10 in = "d";
        #10 in = " ";
        #10 in = "e";
        #10 in = "n";
        #10 in = "d";
        #10 in = " ";
        #5 reset = 1;
        #5 reset = 0;
        #10 in = " ";
        #10 in = "E";
        #10 in = "n";
        #10 in = "d";
        #10 in = " ";
        #10 in = "b";
        #10 in = "E";
        #10 in = "G";
        #10 in = "i";
        #10 in = "n";
        #10 in = " ";
        #10 in = "E";
        #10 in = "n";
        #10 in = "d";
        #10 in = " ";
        #10 in = "E";
        #10 in = "n";
        #10 in = "D";
        #10 in = "E";
        #10 in = " ";
        #10 in = "E";
        #10 in = "n";
        #10 in = "D";
        #10 in = "E";
        #10 in = "n";
        #10 in = "D";
	end
    initial begin
        #500 $finish;
    end
    always #5 clk = ~clk;
endmodule

