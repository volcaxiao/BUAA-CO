`timescale 1ns / 1ps

////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer:
//
// Create Date:   15:11:00 10/06/2022
// Design Name:   gray
// Module Name:   /media/shared/p1/4_gray/gray/gray_tb.v
// Project Name:  gray
// Target Device:  
// Tool versions:  
// Description: 
//
// Verilog Test Fixture created by ISE for module: gray
//
// Dependencies:
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
////////////////////////////////////////////////////////////////////////////////

module gray_tb;

	// Inputs
	reg Clk;
	reg Reset;
	reg En;

	// Outputs
	wire [2:0] Output;
	wire Overflow;

	// Instantiate the Unit Under Test (UUT)
	gray uut (
		.Clk(Clk), 
		.Reset(Reset), 
		.En(En), 
		.Output(Output), 
		.Overflow(Overflow)
	);

	initial begin
		// Initialize Inputs
		Clk = 0;
		Reset = 0;
		En = 0;
		// Wait 100 ns for global reset to finish
        #100
		// Add stimulus here
        En = 1;
        #20 Reset = 1'b1;
        #10 Reset = 1'b0;
        #100 Reset = 1'b1;
        #10 Reset = 1'b0;
	end
   
always #5 Clk = ~Clk;
initial begin
    #300 $finish;
end
endmodule

